/*
 *  GPL-3.0
 *  Copyright (C) 2021  ZaViBiS
 */
module version

pub const version = 0.1
pub const version_url = 'https://raw.githubusercontent.com/ZaViBiS/Percentage-difference/master/version/version.txt'
